module EXC_add  (
    output  wire     [31:0]  Address
);

    assign Address = 32'h88;
    
endmodule